`timescale 1ns / 1ps

module Park_Transform(
    input signed [15:0] i_alpha, i_beta,
    input signed [15:0] sin_theta, cos_theta,
    output reg signed [15:0] i_d, i_q
    );
    
    
    
endmodule
